`default_nettype none
`timescale 1ns/1ps

/*
this testbench just instantiates the module and makes some convenient wires
that can be driven / tested by the cocotb test.py
*/

module tb (
    // testbench is controlled by test.py
    input clk,
    input rst,
    input start, 
    input stop,
    output uart_tx
   );

    // this part dumps the trace to a vcd file that can be viewed with GTKWave
    initial begin
        $dumpfile ("tb.vcd");
        $dumpvars (0, tb);
        #10000;
    end

    // wire up the inputs and outputs
    wire [7:0] inputs = {6'b0,stop, start, rst, clk};
    wire [7:0] outputs;
    assign uart_tx = outputs[0];

    // instantiate the DUT
    Naviss_top top(
        .io_in  (inputs),
        .io_out (outputs)
        );

endmodule
